module counter ( gnd, vdd, enable, clk, reset, out);

input gnd, vdd;
input enable;
input clk;
input reset;
output [7:0] out;

	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(_28__0_), .Y(_1_) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_2_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_3_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(_28__0_), .C(_3_), .Y(_4_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_4_), .Y(_0__0_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(_28__0_), .C(_28__1_), .Y(_5_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_6_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_28__1_), .B(_2_), .C(_3_), .Y(_7_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_7_), .Y(_0__1_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_28__2_), .Y(_8_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_28__1_), .B(_28__2_), .Y(_9_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_9_), .C(_3_), .Y(_10_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_5_), .C(_10_), .Y(_0__2_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_9_), .Y(_11_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_28__3_), .B(_11_), .C(_3_), .Y(_12_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_28__3_), .B(_11_), .C(_12_), .Y(_0__3_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_13_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_28__3_), .B(_28__4_), .Y(_14_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_13_), .Y(_15_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_28__3_), .C(_28__4_), .Y(_16_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_16_), .C(_15_), .Y(_0__4_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_28__5_), .Y(_17_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_13_), .C(_17_), .Y(_18_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_28__3_), .B(_28__4_), .C(_28__5_), .Y(_19_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_20_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_20_), .Y(_21_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_21_), .Y(_22_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_18_), .Y(_0__5_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_28__6_), .B(_21_), .C(_3_), .Y(_23_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_28__6_), .B(_21_), .C(_23_), .Y(_0__6_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_28__6_), .B(_28__7_), .C(_21_), .Y(_24_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_28__7_), .Y(_25_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_28__6_), .B(_20_), .C(_11_), .Y(_26_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_25_), .C(reset), .Y(_27_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_24_), .Y(_0__7_) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_28__0_), .Y(out[0]) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_28__1_), .Y(out[1]) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_28__2_), .Y(out[2]) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_28__3_), .Y(out[3]) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_28__4_), .Y(out[4]) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_28__5_), .Y(out[5]) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_28__6_), .Y(out[6]) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_28__7_), .Y(out[7]) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__0_), .Q(_28__0_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__1_), .Q(_28__1_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__2_), .Q(_28__2_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__3_), .Q(_28__3_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__4_), .Q(_28__4_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__5_), .Q(_28__5_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__6_), .Q(_28__6_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0__7_), .Q(_28__7_) );
endmodule
